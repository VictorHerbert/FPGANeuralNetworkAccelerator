module act_function #(parameter DEPTH)(
    input [DEPTH-1: 0] x,
    output [DEPTH-1: 0] y
);

    assign y = x;
    
endmodule